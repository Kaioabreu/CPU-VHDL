----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create 

